module testMain();
	reg [31:0] a ; // a = 40 ;
	//$display("Decimal value a is: '%d'", a);
endmodule
